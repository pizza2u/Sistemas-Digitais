-- ENGENHARIA ELÉTRICA - IFPB
-- SISTEMAS DIGITAIS 2020.2
-- MINI-PROJETO DA SEMANA 11 (01/05/2021)
-- "PROBLEM 8.3 FROM CIRCUIT DESIGN WITH VHDL"


LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY TESTBENCH IS
END TESTBENCH;

ARCHITECTURE TEST OF TESTBENCH IS

COMPONENT GERADOR IS

PORT(CLK,STOP,GO: IN STD_LOGIC;
     UP,DOWN: OUT STD_LOGIC);

END COMPONENT;

SIGNAL CLOCK,STOP, GO: STD_LOGIC:='0';
SIGNAL UP, DOWN: STD_LOGIC:='0';

BEGIN

DUT: GERADOR PORT MAP(CLOCK,STOP,GO,UP,DOWN);

STOP <= '1', '0' AFTER 30 MS;
             
GO <= '0',
      '1' AFTER 90 MS,
      '0' AFTER 120 MS;
      
	PROCESS
   		
        BEGIN
      	
        FOR I IN 0 TO 70 LOOP
	  	   CLOCK <= '0';
	  	   WAIT FOR 1 MS;
	  	   CLOCK <= '1';
	  	   WAIT FOR 1 MS;
      	END LOOP;
    	
        WAIT;

	END PROCESS; 
 
END TEST;
